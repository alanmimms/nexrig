* Three-Tank BPF Simulation - Simplified
* BAND_NAME

.include BAND_FILE

* Input source
Vin in 0 AC 1

* Input transformer (L1 serves as tank inductor AND transformer secondary)
Lpri in 0 {Ltank/4}
L1 tank1 0 {Ltank}
K1 Lpri L1 0.98

* Tank 1 capacitor
C1 tank1 0 {CtankEnd}

* Coupling C12
C12 tank1 tank2 {Ccouple}

* Tank 2
L2 tank2 0 {Ltank}
C2 tank2 0 {CtankMid}

* Coupling C23
C23 tank2 tank3 {Ccouple}

* Tank 3 - L3 is the transformer secondary
C3 tank3 0 {CtankEnd}

* Output transformer (L3 serves as tank inductor AND transformer secondary)
L3 tank3 0 {Ltank}
Lpri_out out 0 {Ltank/4}
K2 L3 Lpri_out 0.98

* Load
Rload out 0 50

.control
ac dec 100 1MEG 50MEG
set wr_vecnames
set wr_singlescale
wrdata OUTPUT_FILE frequency db(v(out)/v(in))
quit
.endc

.end