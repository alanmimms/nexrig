.title KiCad schematic
.include "/home/alan/ham/usb-ssb-txcvr/spice-models/rn242sm_SPICE.lib"
.save all
.probe alli
.probe p(R7727)
.probe p(R7730)
.probe p(C7831)
.probe p(R7749)
.probe p(I7701)
.probe p(R7748)
.probe p(V7705)
.probe p(L7755)
.probe p(V7704)
.probe p(R7731)
.probe p(V7701)
.probe p(R7733)
.probe p(V7702)
.probe p(C7855)
.probe p(C7856)
.probe p(L7766)
.probe p(L7767)
.probe p(C7851)
.probe p(C7854)
.probe p(L7765)
.probe p(C7850)
.probe p(C7853)
.probe p(C7852)
.probe p(C7849)
.probe p(L7768)
.probe p(D7719)
.probe p(C7859)
.probe p(C7858)
.probe p(C7857)
.probe p(L7769)
.probe p(R7737)
.probe p(D7718)
.probe p(C7846)
.probe p(C7848)
.probe p(L7763)
.probe p(C7847)
.probe p(L7764)
.probe p(R7736)
.probe p(C7883)
.probe p(C7884)
.probe p(L7780)
.probe p(L7781)
.probe p(C7879)
.probe p(C7882)
.probe p(L7779)
.probe p(C7878)
.probe p(C7881)
.probe p(C7880)
.probe p(C7877)
.probe p(L7782)
.probe p(D7723)
.probe p(C7887)
.probe p(C7886)
.probe p(C7885)
.probe p(L7783)
.probe p(R7741)
.probe p(D7722)
.probe p(C7874)
.probe p(C7876)
.probe p(L7777)
.probe p(C7875)
.probe p(L7778)
.probe p(R7740)
.probe p(L2)
.probe p(C2)
.probe p(C4)
.probe p(C3)
.probe p(R7751)
.probe p(L3)
.probe p(C5)
.probe p(L1)
.probe p(V7706)
.probe p(R7750)
.probe p(C7941)
.probe p(L7809)
.probe p(C7935)
.probe p(C7943)
.probe p(C1)
.param Ccouple = 47.8p
.param CtankMid = 68.8p
.param CtankEnd = 116.6p
.ac dec 5000 8Meg 22Meg
R7727 /frontend-sim/Rx_Front_End/RxRFFiltered GND 50
R7730 /frontend-sim/testOut GND 1Meg
C7831 /frontend-sim/testOut GND 385.5p
R7749 /frontend-sim/vLadderOut GND 50
I7701 /frontend-sim/testOut GND DC 0 SIN( 0 1 1k 0 0 0 ) AC 1  
R7748 Net-_R7748-Pad1_ /frontend-sim/test/ladderIn 50
V7705 Net-_R7748-Pad1_ GND DC 0 SIN( 0 1 1k 0 0 0 ) AC 1  
L7755 /frontend-sim/testOut GND 4.7u
V7704 Net-_R7731-Pad1_ GND DC 0 SIN( 0 1 1k 0 0 0 ) AC 1  
R7731 Net-_R7731-Pad1_ /frontend-sim/Rx_Front_End/AntRx 50
V7701 +3.3V GND DC 3.3 
R7733 GND /frontend-sim/RxRFout 50
V7702 +10V GND DC 10 
C7855 Net-_C7854-Pad2_ Net-_C7855-Pad2_ 510p
C7856 Net-_C7855-Pad2_ GND 1500p
L7766 Net-_C7851-Pad2_ GND 4.7u
L7767 Net-_C7854-Pad2_ GND 4.7u
C7851 Net-_C7847-Pad1_ Net-_C7851-Pad2_ 47p
C7854 Net-_C7851-Pad2_ Net-_C7854-Pad2_ 47p
L7765 Net-_C7847-Pad1_ GND 4.7u
C7850 Net-_C7847-Pad1_ Net-_C7847-Pad2_ 1f
C7853 Net-_C7851-Pad2_ GND 30.156p
C7852 Net-_C7851-Pad2_ GND 330p
C7849 Net-_C7847-Pad2_ GND 100p
L7768 GND Net-_C7855-Pad2_ 470u
D7719 Net-_C7855-Pad2_ Net-_C7859-Pad1_ DRN242SM
C7859 Net-_C7859-Pad1_ /frontend-sim/Rx_Front_End/RxRFFiltered 0.1u
C7858 Net-_C7855-Pad2_ GND 100p
C7857 Net-_C7854-Pad2_ Net-_C7855-Pad2_ 1f
L7769 Net-_L7769-Pad1_ GND 470u
R7737 Net-_L7769-Pad1_ Net-_C7859-Pad1_ 680
D7718 Net-_C7846-Pad2_ Net-_C7847-Pad2_ DRN242SM
C7846 /frontend-sim/Rx_Front_End/AntRx Net-_C7846-Pad2_ 0.1u
C7848 Net-_C7847-Pad2_ GND 1500p
L7763 GND Net-_C7846-Pad2_ 470u
C7847 Net-_C7847-Pad1_ Net-_C7847-Pad2_ 510p
L7764 Net-_L7764-Pad1_ GND 470u
R7736 Net-_L7764-Pad1_ Net-_C7847-Pad2_ 680
C7883 Net-_C7882-Pad2_ Net-_C7883-Pad2_ 150p
C7884 Net-_C7883-Pad2_ GND 220p
L7780 Net-_C7879-Pad2_ GND 1u
L7781 Net-_C7882-Pad2_ GND 1u
C7879 Net-_C7875-Pad1_ Net-_C7879-Pad2_ 25p
C7882 Net-_C7879-Pad2_ Net-_C7882-Pad2_ 25p
L7779 Net-_C7875-Pad1_ GND 1u
C7878 Net-_C7875-Pad1_ Net-_C7875-Pad2_ 1f
C7881 Net-_C7879-Pad2_ GND 30.156p
C7880 Net-_C7879-Pad2_ GND 82p
C7877 Net-_C7875-Pad2_ GND 47p
L7782 +3.3V Net-_C7883-Pad2_ 470u
D7723 Net-_C7883-Pad2_ Net-_C7887-Pad1_ DRN242SM
C7887 Net-_C7887-Pad1_ /frontend-sim/Rx_Front_End/RxRFFiltered 0.1u
C7886 Net-_C7883-Pad2_ GND 47p
C7885 Net-_C7882-Pad2_ Net-_C7883-Pad2_ 1f
L7783 Net-_L7783-Pad1_ GND 470u
R7741 Net-_L7783-Pad1_ Net-_C7887-Pad1_ 680
D7722 Net-_C7874-Pad2_ Net-_C7875-Pad2_ DRN242SM
C7874 /frontend-sim/Rx_Front_End/AntRx Net-_C7874-Pad2_ 0.1u
C7876 Net-_C7875-Pad2_ GND 220p
L7777 +3.3V Net-_C7874-Pad2_ 470u
C7875 Net-_C7875-Pad1_ Net-_C7875-Pad2_ 150p
L7778 Net-_L7778-Pad1_ GND 470u
R7740 Net-_L7778-Pad1_ Net-_C7875-Pad2_ 680
L2 Net-_C2-Pad2_ GND 617n
C2 Net-_C1-Pad1_ Net-_C2-Pad2_ {Ccouple}
C4 Net-_C2-Pad2_ /frontend-sim/test/vACOut {Ccouple}
C3 Net-_C2-Pad2_ GND {CtankMid}
R7751 /frontend-sim/test/vACOut GND 200
L3 /frontend-sim/test/vACOut GND 617n
C5 /frontend-sim/test/vACOut GND {CtankEnd}
L1 Net-_C1-Pad1_ GND 617n
V7706 Net-_R7750-Pad2_ GND DC 0 SIN( 0 1 1k 0 0 0 ) AC 1  
R7750 Net-_C1-Pad1_ Net-_R7750-Pad2_ 200
C7941 Net-_C7941-Pad1_ /frontend-sim/vLadderOut 126.084p
L7809 /frontend-sim/test/ladderIn Net-_C7941-Pad1_ 1u
C7935 /frontend-sim/test/ladderIn GND 9381.96p
C7943 /frontend-sim/vLadderOut GND 9381.96p
C1 Net-_C1-Pad1_ GND {CtankEnd}
.end

.control
set noaskquit

let Cvals = vector(80p, 90p, 100p, 110p, 120p, 130p, 140p, 150p)
foreach c $&Cvals
    alterparam CtankEnd = c
    run
end
.endc

