* Simple 3rd-order LPF test - should show steep rolloff
* Using Band 1 values

.param L1=6533n
.param C1=243p  
.param L2=6533n

V1 in 0 AC 1 0
Rs in n1 50

* Simple 3rd-order LPF (no transformers)
L1 n1 n2 {L1}
C1 n2 0 {C1}
L2 n2 n3 {L2}
Rload n3 0 200

.ac dec 100 100k 100meg
.control
run
print frequency vdb(n3)
.endc
.end