* Working 40m 3-Pole BPF - CORRECT Topology
* Transformer-coupled three-tank design

.param L=106103n
.param C_main=6p
.param C_tap=19p
.param C_couple=0p

* === SOURCE ===
V1 in 0 AC 1 0
Rs in n1 50

* === 3-TANK BANDPASS FILTER ===
* Tank 1: Input tank with tapped capacitor for 50Ω matching
L1 n2 n3 {L}
C1_main n3 0 {C_main}
C1_tap n1 n2 {C_tap}

* Tank 2: Center tank (parallel resonant)
L2 n4 n5 {L}
C2 n5 0 {C_main}

* Tank 3: Output tank with tapped capacitor for 50Ω matching  
L3 n6 n7 {L}
C3_main n7 0 {C_main}
C3_tap n6 n8 {C_tap}

* Coupling between tanks
C12 n3 n4 {C_couple}  ; Tank 1 to Tank 2
C23 n5 n6 {C_couple}  ; Tank 2 to Tank 3

* === LOAD ===
RL n8 0 50

* === ANALYSIS ===
.ac dec 100 1meg 100meg
.control
run
print frequency vdb(n8)
.endc
.end
